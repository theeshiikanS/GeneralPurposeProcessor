library verilog;
use verilog.vl_types.all;
entity ALU2Schematic_vlg_vec_tst is
end ALU2Schematic_vlg_vec_tst;
